`timescale 1ns/1ps
`celldefine
//
// I_FAB simulation model
// Marker Buffer for periphery to fabric transition
//
// Copyright (c) 2024 Rapid Silicon, Inc.  All rights reserved.
//

module I_FAB (
  input I, // Input
  output O // Output
);

assign O = I ;


endmodule
`endcelldefine
