`timescale 1ns/1ps
`celldefine
//
// O_FAB simulation model
// Marker Buffer for fabric to pheriphery transition 
//
// Copyright (c) 2024 Rapid Silicon, Inc.  All rights reserved.
//

module O_FAB (
  input I, // Input
  output O // Output
);

   assign O = I ;

endmodule
`endcelldefine
